module iQueue(
    input i_drive,
    input[7*0] i_cutPostion_8,
    input[32*10-1:0] i_alignedInstructionTable,
    output 
);

    reg[31:0] q[15:0];

    
endmodule